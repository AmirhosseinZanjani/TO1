magic
tech sky130A
magscale 1 2
timestamp 1696943305
<< nwell >>
rect -13652 8716 -13602 8762
rect -16204 7948 -16098 7982
rect -14646 7954 -14408 7982
rect -14664 7898 -14636 7950
rect -16240 7758 -16194 7846
rect -14664 7758 -14626 7844
<< pwell >>
rect -16974 7446 -12742 7466
rect -17838 7436 -12742 7446
rect -17838 7420 -12454 7436
rect -17838 6744 -17830 7420
rect -12514 7282 -12508 7284
rect -17690 6744 -16748 6842
rect -15148 6768 -15144 6892
rect -15144 6758 -15124 6764
rect -13428 6744 -13394 6842
rect -12850 6808 -12816 6944
rect -12476 6744 -12454 7420
rect -17838 6706 -12454 6744
rect -16736 6682 -12454 6706
rect -16736 6640 -13508 6682
rect -16760 6572 -13508 6640
<< psubdiff >>
rect -16974 7446 -12742 7464
rect -17838 7436 -12742 7446
rect -17838 7420 -12500 7436
rect -17838 6888 -17830 7420
<< locali >>
rect -18008 8944 -12356 9382
rect -18008 8942 -13660 8944
rect -18008 8892 -16750 8942
rect -18008 7898 -17862 8892
rect -16688 8924 -13660 8942
rect -16688 8892 -15206 8924
rect -17728 8786 -16756 8824
rect -16548 8788 -16504 8892
rect -15144 8892 -13660 8924
rect -13598 8892 -12356 8944
rect -16432 8788 -15492 8822
rect -14792 8788 -13914 8822
rect -13840 8786 -13796 8892
rect -12496 8848 -12358 8892
rect -13526 8788 -12610 8826
rect -12500 8762 -12358 8848
rect -12496 8574 -12358 8762
rect -18006 7792 -17862 7898
rect -16394 7855 -16282 7890
rect -16082 7855 -15814 7890
rect -15618 7855 -15460 7890
rect -14890 7860 -13920 7893
rect -12498 7860 -12358 8574
rect -14890 7853 -14020 7860
rect -18006 7756 -16248 7792
rect -16186 7756 -15708 7792
rect -15646 7758 -14674 7792
rect -14612 7758 -14176 7792
rect -15646 7756 -14176 7758
rect -12496 7792 -12358 7860
rect -14114 7756 -12358 7792
rect -18006 7664 -12358 7756
rect -18006 7660 -17862 7664
rect -17838 7436 -12742 7446
rect -17838 7420 -12454 7436
rect -17838 6744 -17830 7420
rect -16378 7318 -15702 7352
rect -15646 7318 -14671 7353
rect -14606 7320 -13896 7358
rect -12476 7290 -12454 7420
rect -17494 6842 -17460 6946
rect -12850 6842 -12816 6944
rect -12594 6882 -12570 7128
rect -12480 6862 -12454 7290
rect -17690 6744 -16748 6842
rect -16420 6798 -15710 6836
rect -15644 6804 -15470 6842
rect -14800 6804 -14668 6842
rect -14606 6802 -13896 6840
rect -13578 6808 -12620 6842
rect -17838 6726 -15172 6744
rect -17838 6710 -15308 6726
rect -17838 6706 -16002 6710
rect -13574 6744 -12620 6808
rect -12476 6744 -12454 6862
rect -15138 6726 -12454 6744
rect -13820 6724 -12454 6726
<< viali >>
rect -16750 8890 -16688 8942
rect -15206 8872 -15144 8924
rect -13660 8892 -13598 8944
rect -16248 7756 -16186 7808
rect -15708 7756 -15646 7808
rect -14674 7758 -14612 7810
rect -14176 7756 -14114 7808
rect -15172 6706 -15138 6746
<< metal1 >>
rect -16760 8942 -16678 8954
rect -16760 8890 -16750 8942
rect -16688 8890 -16678 8942
rect -13670 8944 -13588 8956
rect -16760 8878 -16678 8890
rect -15218 8924 -15130 8940
rect -15218 8872 -15206 8924
rect -15144 8872 -15130 8924
rect -13670 8892 -13660 8944
rect -13598 8892 -13588 8944
rect -13670 8880 -13588 8892
rect -15218 8860 -15130 8872
rect -17434 8788 -17424 8856
rect -17274 8788 -17264 8856
rect -16130 8784 -16120 8852
rect -15970 8784 -15960 8852
rect -15352 8788 -15342 8842
rect -15290 8788 -15280 8842
rect -15090 8788 -15080 8842
rect -15028 8788 -15018 8842
rect -14348 8790 -14338 8858
rect -14188 8790 -14178 8858
rect -13040 8784 -13030 8852
rect -12880 8784 -12870 8852
rect -15982 8718 -15972 8720
rect -17788 8662 -17778 8716
rect -17726 8662 -17716 8716
rect -17274 8662 -17264 8716
rect -17212 8662 -17202 8716
rect -16766 8662 -16756 8716
rect -16704 8662 -16694 8716
rect -16502 8632 -16492 8718
rect -16430 8632 -16420 8718
rect -15986 8630 -15976 8718
rect -15914 8632 -15904 8720
rect -15918 8630 -15908 8632
rect -15478 8628 -15468 8714
rect -15406 8628 -15396 8714
rect -15210 8696 -15200 8750
rect -15148 8696 -15138 8750
rect -14952 8628 -14942 8714
rect -14880 8628 -14870 8714
rect -14440 8624 -14430 8712
rect -14372 8624 -14362 8712
rect -13924 8624 -13914 8712
rect -13856 8624 -13846 8712
rect -13660 8664 -13650 8718
rect -13598 8664 -13588 8718
rect -13142 8664 -13132 8718
rect -13080 8664 -13070 8718
rect -12628 8664 -12618 8718
rect -12566 8664 -12556 8718
rect -17522 8228 -17512 8314
rect -17450 8228 -17440 8314
rect -17014 8218 -17004 8304
rect -16942 8218 -16932 8304
rect -13396 8230 -13386 8316
rect -13324 8230 -13314 8316
rect -12890 8218 -12880 8304
rect -12818 8218 -12808 8304
rect -16258 7946 -16248 7998
rect -16186 7946 -16176 7998
rect -15734 7946 -15724 7998
rect -15662 7946 -15652 7998
rect -14686 7944 -14682 8034
rect -14674 7938 -14664 7990
rect -14602 7938 -14592 7990
rect -14186 7938 -14176 7990
rect -14114 7938 -14104 7990
rect -15580 7826 -15570 7896
rect -15454 7826 -15444 7896
rect -14884 7826 -14874 7896
rect -14758 7826 -14748 7896
rect -16260 7808 -16174 7820
rect -16260 7756 -16248 7808
rect -16186 7756 -16174 7808
rect -16260 7744 -16174 7756
rect -15724 7808 -15636 7820
rect -15724 7756 -15708 7808
rect -15646 7756 -15636 7808
rect -15724 7744 -15636 7756
rect -14684 7810 -14602 7822
rect -14684 7758 -14674 7810
rect -14612 7758 -14602 7810
rect -14684 7746 -14602 7758
rect -14186 7808 -14104 7820
rect -14186 7756 -14176 7808
rect -14114 7756 -14104 7808
rect -14186 7744 -14104 7756
rect -15592 7296 -15582 7374
rect -15484 7296 -15474 7374
rect -14832 7296 -14822 7374
rect -14724 7296 -14714 7374
rect -16222 7208 -16212 7277
rect -16158 7208 -16148 7277
rect -15712 7207 -15702 7276
rect -15648 7207 -15638 7276
rect -15192 7256 -15183 7277
rect -15193 7208 -15183 7256
rect -15129 7252 -15120 7277
rect -14674 7252 -14667 7276
rect -15129 7208 -15119 7252
rect -14677 7207 -14667 7252
rect -14613 7207 -14603 7276
rect -14160 7212 -14150 7281
rect -14096 7212 -14086 7281
rect -17768 7036 -17758 7105
rect -17704 7036 -17694 7105
rect -17252 7056 -17242 7107
rect -17248 7038 -17242 7056
rect -17188 7038 -17178 7107
rect -16734 7064 -16724 7105
rect -16732 7036 -16724 7064
rect -16670 7036 -16660 7105
rect -16473 7036 -16463 7105
rect -16409 7036 -16399 7105
rect -15966 7034 -15956 7103
rect -15902 7034 -15892 7103
rect -14415 7039 -14405 7108
rect -14351 7039 -14341 7108
rect -13907 7032 -13897 7101
rect -13843 7032 -13833 7101
rect -13638 7038 -13628 7107
rect -13574 7038 -13564 7107
rect -13122 7040 -13112 7109
rect -13058 7040 -13048 7109
rect -12610 7036 -12600 7105
rect -12546 7036 -12536 7105
rect -17512 6886 -17502 6938
rect -17440 6886 -17430 6938
rect -17002 6886 -16992 6938
rect -16930 6886 -16920 6938
rect -15444 6886 -15434 6938
rect -15372 6886 -15362 6938
rect -14932 6886 -14922 6938
rect -14860 6886 -14850 6938
rect -13384 6890 -13374 6942
rect -13312 6890 -13302 6942
rect -12866 6890 -12856 6942
rect -12794 6890 -12786 6942
rect -16610 6750 -16600 6844
rect -16488 6750 -16478 6844
rect -13786 6792 -13776 6870
rect -13700 6792 -13690 6870
rect -13578 6808 -13498 6842
rect -15196 6706 -15186 6758
rect -15124 6706 -15114 6758
rect -15196 6696 -15114 6706
<< via1 >>
rect -16750 8890 -16688 8942
rect -15206 8872 -15144 8924
rect -13660 8892 -13598 8944
rect -17424 8788 -17274 8856
rect -16120 8784 -15970 8852
rect -15342 8788 -15290 8842
rect -15080 8788 -15028 8842
rect -14338 8790 -14188 8858
rect -13030 8784 -12880 8852
rect -15972 8718 -15914 8720
rect -17778 8662 -17726 8716
rect -17264 8662 -17212 8716
rect -16756 8662 -16704 8716
rect -16492 8632 -16430 8718
rect -15976 8632 -15914 8718
rect -15976 8630 -15918 8632
rect -15468 8628 -15406 8714
rect -15200 8696 -15148 8750
rect -14942 8628 -14880 8714
rect -14430 8624 -14372 8712
rect -13914 8624 -13856 8712
rect -13650 8664 -13598 8718
rect -13132 8664 -13080 8718
rect -12618 8664 -12566 8718
rect -17512 8228 -17450 8314
rect -17004 8218 -16942 8304
rect -13386 8230 -13324 8316
rect -12880 8218 -12818 8304
rect -16248 7946 -16186 7998
rect -15724 7946 -15662 7998
rect -14664 7938 -14602 7990
rect -14176 7938 -14114 7990
rect -15570 7826 -15454 7896
rect -14874 7826 -14758 7896
rect -16248 7756 -16186 7808
rect -15708 7756 -15646 7808
rect -14674 7758 -14612 7810
rect -14176 7756 -14114 7808
rect -15582 7296 -15484 7374
rect -14822 7296 -14724 7374
rect -16212 7208 -16158 7277
rect -15702 7207 -15648 7276
rect -15183 7208 -15129 7277
rect -14667 7207 -14613 7276
rect -14150 7212 -14096 7281
rect -17758 7036 -17704 7105
rect -17242 7038 -17188 7107
rect -16724 7036 -16670 7105
rect -16463 7036 -16409 7105
rect -15956 7034 -15902 7103
rect -14405 7039 -14351 7108
rect -13897 7032 -13843 7101
rect -13628 7038 -13574 7107
rect -13112 7040 -13058 7109
rect -12600 7036 -12546 7105
rect -17502 6886 -17440 6938
rect -16992 6886 -16930 6938
rect -15434 6886 -15372 6938
rect -14922 6886 -14860 6938
rect -13374 6890 -13312 6942
rect -12856 6890 -12794 6942
rect -16600 6750 -16488 6844
rect -13776 6792 -13700 6870
rect -15186 6746 -15124 6758
rect -15186 6706 -15172 6746
rect -15172 6706 -15138 6746
rect -15138 6706 -15124 6746
<< metal2 >>
rect -17386 9132 -17302 9142
rect -17386 9052 -17302 9062
rect -16072 9132 -15988 9142
rect -16072 9052 -15988 9062
rect -14286 9132 -14202 9142
rect -14286 9052 -14202 9062
rect -12988 9132 -12904 9142
rect -12988 9052 -12904 9062
rect -17386 8880 -17338 9052
rect -16750 8942 -16688 8952
rect -16750 8880 -16688 8890
rect -17386 8868 -17306 8880
rect -17416 8866 -17280 8868
rect -17424 8856 -17274 8866
rect -17424 8778 -17274 8788
rect -16740 8730 -16706 8880
rect -16072 8868 -16012 9052
rect -15452 8974 -15012 9016
rect -16072 8864 -15974 8868
rect -16110 8862 -15974 8864
rect -16120 8852 -15970 8862
rect -16120 8774 -15970 8784
rect -16740 8726 -16704 8730
rect -15972 8728 -15914 8730
rect -16492 8726 -16430 8728
rect -17778 8716 -17726 8726
rect -17264 8716 -17212 8726
rect -16756 8716 -16704 8726
rect -17726 8662 -17264 8716
rect -17212 8662 -16756 8716
rect -17778 8652 -17726 8662
rect -17264 8652 -17212 8662
rect -16756 8652 -16704 8662
rect -16494 8718 -16430 8726
rect -15976 8720 -15914 8728
rect -15452 8724 -15416 8974
rect -15206 8924 -15144 8934
rect -15362 8856 -15264 8866
rect -15206 8862 -15144 8872
rect -15362 8768 -15264 8778
rect -15198 8760 -15152 8862
rect -15090 8842 -15012 8974
rect -14286 8866 -14218 9052
rect -13660 8944 -13598 8954
rect -13660 8882 -13598 8892
rect -15090 8790 -15080 8842
rect -15028 8790 -15012 8842
rect -14338 8858 -14188 8866
rect -15080 8778 -15028 8788
rect -14338 8780 -14188 8790
rect -15200 8750 -15148 8760
rect -15976 8718 -15972 8720
rect -15468 8718 -15406 8724
rect -16494 8716 -16492 8718
rect -16430 8632 -15976 8718
rect -15914 8714 -15406 8718
rect -15914 8632 -15468 8714
rect -16434 8630 -15976 8632
rect -15918 8630 -15468 8632
rect -16434 8628 -15468 8630
rect -13652 8728 -13602 8882
rect -12980 8862 -12906 9052
rect -13030 8852 -12880 8862
rect -13030 8774 -12880 8784
rect -15200 8686 -15148 8696
rect -14942 8714 -14880 8724
rect -14430 8714 -14372 8722
rect -13914 8714 -13856 8722
rect -13652 8718 -13598 8728
rect -13652 8716 -13650 8718
rect -16434 8622 -16430 8628
rect -15976 8622 -15914 8628
rect -15494 8626 -15406 8628
rect -15976 8620 -15918 8622
rect -16494 8610 -16434 8620
rect -15468 8618 -15406 8626
rect -14880 8712 -13856 8714
rect -14880 8628 -14430 8712
rect -14942 8624 -14430 8628
rect -14372 8704 -13914 8712
rect -14372 8624 -13920 8704
rect -13132 8718 -13080 8728
rect -13598 8664 -13132 8716
rect -12618 8718 -12566 8728
rect -13080 8664 -12618 8716
rect -13650 8662 -12566 8664
rect -13650 8654 -13598 8662
rect -13132 8654 -13080 8662
rect -12618 8654 -12566 8662
rect -14942 8622 -14780 8624
rect -14942 8618 -14880 8622
rect -14430 8614 -14372 8624
rect -13858 8618 -13856 8624
rect -13920 8614 -13856 8618
rect -13920 8608 -13858 8614
rect -17512 8314 -17450 8324
rect -13386 8316 -13324 8326
rect -17520 8228 -17512 8314
rect -17004 8308 -16942 8314
rect -17450 8304 -16942 8308
rect -17450 8228 -17004 8304
rect -17520 8218 -17004 8228
rect -13392 8230 -13386 8316
rect -13324 8314 -12838 8316
rect -13324 8304 -12818 8314
rect -13324 8230 -12880 8304
rect -13392 8226 -12880 8230
rect -13386 8220 -13324 8226
rect -17520 7632 -17468 8218
rect -17004 8208 -16942 8218
rect -12880 8208 -12818 8218
rect -16248 7998 -16186 8008
rect -15724 7998 -15662 8008
rect -16186 7948 -15724 7982
rect -16248 7936 -16186 7946
rect -14664 7990 -14602 8000
rect -15724 7936 -15662 7946
rect -16240 7818 -16194 7936
rect -15702 7818 -15662 7936
rect -15570 7962 -15454 7972
rect -16248 7808 -16186 7818
rect -16248 7746 -16186 7756
rect -15708 7808 -15646 7818
rect -15570 7816 -15454 7826
rect -14874 7970 -14758 7980
rect -14874 7816 -14758 7826
rect -14176 7990 -14114 8000
rect -14602 7954 -14176 7982
rect -14664 7928 -14602 7938
rect -14176 7928 -14114 7938
rect -14664 7848 -14624 7928
rect -14664 7820 -14626 7848
rect -15708 7746 -15646 7756
rect -14674 7810 -14612 7820
rect -14170 7818 -14134 7928
rect -14674 7748 -14612 7758
rect -14176 7808 -14114 7818
rect -14176 7746 -14114 7756
rect -12878 7636 -12826 8208
rect -17526 7580 -16416 7632
rect -13894 7588 -12828 7636
rect -17520 7578 -17468 7580
rect -16732 7372 -16672 7382
rect -16732 7266 -16672 7276
rect -17758 7112 -17704 7115
rect -17242 7112 -17188 7117
rect -16726 7115 -16682 7266
rect -16462 7122 -16418 7580
rect -15582 7374 -15484 7384
rect -16212 7277 -16158 7287
rect -15582 7286 -15484 7296
rect -14822 7374 -14724 7384
rect -16227 7219 -16212 7274
rect -15702 7276 -15648 7286
rect -16158 7219 -15702 7274
rect -16212 7198 -16158 7208
rect -15183 7277 -15129 7287
rect -14822 7286 -14724 7296
rect -15648 7256 -15638 7274
rect -15192 7256 -15183 7273
rect -15648 7220 -15183 7256
rect -15648 7219 -15624 7220
rect -15702 7197 -15648 7207
rect -14667 7276 -14613 7286
rect -15129 7252 -15120 7273
rect -14674 7252 -14667 7273
rect -15129 7220 -14667 7252
rect -15183 7198 -15129 7208
rect -14150 7281 -14096 7291
rect -14613 7220 -14150 7273
rect -14667 7197 -14613 7207
rect -14096 7220 -14077 7273
rect -14150 7202 -14096 7212
rect -13894 7122 -13852 7588
rect -12878 7586 -12828 7588
rect -13642 7370 -13582 7380
rect -13582 7274 -13580 7279
rect -13642 7264 -13580 7274
rect -13624 7140 -13580 7264
rect -13628 7130 -13568 7140
rect -16726 7112 -16670 7115
rect -17758 7107 -16670 7112
rect -17758 7105 -17242 7107
rect -17704 7056 -17242 7105
rect -17704 7036 -17692 7056
rect -17758 7034 -17692 7036
rect -17248 7038 -17242 7056
rect -17188 7105 -16670 7107
rect -17188 7064 -16724 7105
rect -17188 7038 -17176 7064
rect -17248 7034 -17176 7038
rect -16732 7036 -16724 7064
rect -16732 7034 -16670 7036
rect -17758 7026 -17704 7034
rect -17242 7028 -17188 7034
rect -16724 7026 -16670 7034
rect -16463 7113 -15912 7122
rect -14397 7118 -13846 7122
rect -16463 7105 -15902 7113
rect -16409 7103 -15902 7105
rect -16409 7036 -15956 7103
rect -16463 7034 -15956 7036
rect -17502 6938 -17440 6944
rect -16992 6938 -16930 6944
rect -17440 6924 -17430 6926
rect -17002 6924 -16992 6926
rect -17440 6896 -16992 6924
rect -17440 6892 -17430 6896
rect -17236 6892 -16992 6896
rect -17502 6880 -17440 6886
rect -16992 6880 -16930 6886
rect -16724 6632 -16686 7026
rect -16463 7024 -15902 7034
rect -14405 7111 -13846 7118
rect -14405 7108 -13843 7111
rect -14351 7101 -13843 7108
rect -14351 7039 -13897 7101
rect -14405 7032 -13897 7039
rect -14405 7029 -13843 7032
rect -16463 7022 -15912 7024
rect -14397 7022 -13843 7029
rect -13112 7110 -13058 7119
rect -12600 7110 -12546 7115
rect -13568 7109 -12546 7110
rect -13568 7040 -13112 7109
rect -13058 7105 -12546 7109
rect -13058 7040 -12600 7105
rect -13568 7036 -12600 7040
rect -13568 7034 -12546 7036
rect -13628 7032 -12546 7034
rect -13628 7024 -13568 7032
rect -13112 7030 -13058 7032
rect -12600 7026 -12546 7032
rect -15434 6938 -15372 6944
rect -14922 6938 -14860 6944
rect -15180 6924 -15128 6926
rect -15372 6892 -14922 6924
rect -15434 6880 -15372 6886
rect -16600 6844 -16488 6854
rect -15172 6764 -15144 6892
rect -14922 6880 -14860 6886
rect -13374 6942 -13312 6948
rect -12856 6942 -12794 6948
rect -13312 6896 -12856 6924
rect -13312 6890 -13302 6896
rect -12866 6890 -12856 6896
rect -13374 6884 -13312 6890
rect -12856 6884 -12794 6890
rect -13776 6870 -13700 6880
rect -13820 6792 -13776 6838
rect -13700 6792 -13652 6838
rect -16600 6740 -16488 6750
rect -15186 6758 -15124 6764
rect -15186 6696 -15124 6706
rect -13820 6696 -13652 6792
rect -13818 6632 -13654 6696
rect -16724 6590 -13654 6632
<< via2 >>
rect -17386 9062 -17302 9132
rect -16072 9062 -15988 9132
rect -14286 9062 -14202 9132
rect -12988 9062 -12904 9132
rect -15362 8842 -15264 8856
rect -15362 8788 -15342 8842
rect -15342 8788 -15290 8842
rect -15290 8788 -15264 8842
rect -15362 8778 -15264 8788
rect -16494 8632 -16492 8716
rect -16492 8632 -16434 8716
rect -16494 8620 -16434 8632
rect -14942 8628 -14880 8714
rect -13920 8624 -13914 8704
rect -13914 8624 -13858 8704
rect -13920 8618 -13858 8624
rect -15570 7896 -15454 7962
rect -15570 7852 -15454 7896
rect -14874 7896 -14758 7970
rect -14874 7860 -14758 7896
rect -16732 7276 -16672 7372
rect -15582 7296 -15484 7374
rect -14822 7296 -14724 7374
rect -13642 7274 -13582 7370
rect -13628 7107 -13568 7130
rect -13628 7038 -13574 7107
rect -13574 7038 -13568 7107
rect -13628 7034 -13568 7038
rect -16600 6750 -16488 6844
<< metal3 >>
rect -17396 9132 -17292 9200
rect -17396 9062 -17386 9132
rect -17302 9062 -17292 9132
rect -17396 9056 -17292 9062
rect -16082 9132 -15978 9200
rect -16082 9062 -16072 9132
rect -15988 9062 -15978 9132
rect -16082 9056 -15978 9062
rect -14296 9132 -14192 9202
rect -14296 9062 -14286 9132
rect -14202 9062 -14192 9132
rect -14296 9057 -14192 9062
rect -12998 9132 -12894 9200
rect -12998 9062 -12988 9132
rect -12904 9062 -12894 9132
rect -12998 9056 -12894 9062
rect -15342 8960 -14878 9026
rect -15342 8866 -15264 8960
rect -15362 8861 -15264 8866
rect -15372 8856 -15254 8861
rect -15372 8778 -15362 8856
rect -15264 8778 -15254 8856
rect -15372 8773 -15254 8778
rect -16524 8716 -16416 8724
rect -14944 8719 -14878 8960
rect -16524 8620 -16494 8716
rect -16434 8620 -16416 8716
rect -14952 8714 -14870 8719
rect -14952 8628 -14942 8714
rect -14880 8628 -14870 8714
rect -13908 8709 -13840 8722
rect -14952 8623 -14870 8628
rect -13930 8704 -13840 8709
rect -16524 8420 -16416 8620
rect -13930 8618 -13920 8704
rect -13858 8618 -13840 8704
rect -13930 8613 -13840 8618
rect -16746 8416 -16416 8420
rect -16748 8326 -16416 8416
rect -13908 8420 -13840 8613
rect -13908 8414 -13578 8420
rect -13908 8326 -13562 8414
rect -16748 7372 -16660 8326
rect -15604 7973 -15468 7975
rect -15604 7962 -15444 7973
rect -15604 7892 -15570 7962
rect -15626 7852 -15570 7892
rect -15454 7892 -15444 7962
rect -14884 7970 -14748 7975
rect -14884 7892 -14874 7970
rect -15454 7852 -15440 7892
rect -15626 7742 -15440 7852
rect -14892 7860 -14874 7892
rect -14758 7892 -14748 7970
rect -14758 7860 -14686 7892
rect -14892 7742 -14686 7860
rect -15626 7740 -15490 7742
rect -15626 7716 -15506 7740
rect -15608 7706 -15506 7716
rect -15596 7452 -15506 7706
rect -14786 7570 -14686 7742
rect -14786 7454 -14684 7570
rect -15596 7404 -15440 7452
rect -14892 7410 -14684 7454
rect -14922 7404 -14684 7410
rect -15596 7400 -14684 7404
rect -16748 7276 -16732 7372
rect -16672 7276 -16660 7372
rect -15626 7388 -14684 7400
rect -15626 7374 -14686 7388
rect -13650 7375 -13562 8326
rect -15626 7318 -15582 7374
rect -15592 7296 -15582 7318
rect -15484 7318 -14822 7374
rect -15484 7296 -15474 7318
rect -15592 7291 -15474 7296
rect -14832 7296 -14822 7318
rect -14724 7318 -14686 7374
rect -13652 7370 -13562 7375
rect -14724 7296 -14714 7318
rect -14832 7291 -14714 7296
rect -16748 7266 -16660 7276
rect -13652 7274 -13642 7370
rect -13582 7274 -13562 7370
rect -13652 7272 -13562 7274
rect -13652 7269 -13572 7272
rect -13638 7130 -13558 7135
rect -13638 7034 -13628 7130
rect -13568 7034 -13558 7130
rect -13638 7029 -13558 7034
rect -16610 6844 -16478 6849
rect -16610 6842 -16600 6844
rect -16670 6750 -16600 6842
rect -16488 6750 -16478 6844
rect -16670 6745 -16478 6750
rect -16670 6660 -16490 6745
rect -13638 6660 -13574 7029
rect -16670 6590 -13574 6660
<< via3 >>
rect -17386 9062 -17302 9132
rect -16072 9062 -15988 9132
rect -14286 9062 -14202 9132
rect -12988 9062 -12904 9132
<< metal4 >>
rect -17396 9062 -17386 9200
rect -16082 9062 -16072 9200
rect -17396 9056 -17292 9062
rect -16082 9056 -15978 9062
rect -14202 9060 -14192 9202
rect -12904 9062 -12892 9202
rect -14296 9057 -14192 9060
rect -12998 9056 -12892 9062
<< via4 >>
rect -17386 9132 -17076 9332
rect -17386 9062 -17302 9132
rect -17302 9062 -17076 9132
rect -16072 9132 -15762 9332
rect -16072 9062 -15988 9132
rect -15988 9062 -15762 9132
rect -14512 9132 -14202 9330
rect -14512 9062 -14286 9132
rect -14286 9062 -14202 9132
rect -14512 9060 -14202 9062
rect -13214 9132 -12904 9332
rect -13214 9062 -12988 9132
rect -12988 9062 -12904 9132
<< metal5 >>
rect -17410 9332 -12878 9382
rect -17410 9062 -17386 9332
rect -17076 9062 -16072 9332
rect -15762 9330 -13214 9332
rect -15762 9062 -14512 9330
rect -17410 9060 -14512 9062
rect -14202 9062 -13214 9330
rect -12904 9062 -12878 9332
rect -14202 9060 -12880 9062
rect -17410 9038 -12880 9060
rect -14536 9036 -14178 9038
use sky130_fd_pr__nfet_01v8_5GHK3V  sky130_fd_pr__nfet_01v8_5GHK3V_0
timestamp 1695733796
transform 1 0 -15155 0 1 7080
box -2747 -410 2747 410
use sky130_fd_pr__pfet_01v8_56UW44  sky130_fd_pr__pfet_01v8_56UW44_0
timestamp 1695705298
transform 1 0 -15175 0 1 8341
box -2747 -619 2747 619
<< labels >>
rlabel space -18192 8876 -15224 9302 1 Vdd
rlabel space -18192 6446 -12284 6842 1 Vss
rlabel space -18020 8876 -15224 9216 1 Vdd
rlabel space -18020 6530 -16732 6742 1 Vss
rlabel space -17914 8876 -15224 9216 1 vdd
rlabel space -17914 6530 -16732 6742 1 vss
rlabel space -17914 6530 -16732 6742 1 Vss
rlabel space -17914 8876 -15224 9216 1 Vdd
rlabel metal2 -17526 7580 -16416 7632 1 nodeA1
rlabel metal2 -13894 7588 -12828 7636 1 nodeA2
rlabel space -17708 6740 -17398 6840 1 Vss
rlabel space -16418 7318 -15702 7352 1 InP
rlabel space -17866 6706 -17770 6740 1 Vss
rlabel locali -14606 7320 -13896 7358 1 InN
rlabel metal2 -13568 7032 -13112 7110 1 OP
rlabel space -17188 7034 -16724 7112 1 ON
rlabel metal2 -16158 7219 -15702 7274 1 net1
rlabel space -17886 7854 -17852 8828 1 Vdd
rlabel locali -15646 7318 -14671 7353 1 Clk
rlabel metal2 -15198 8750 -15152 8872 1 vdd
rlabel metal3 -13650 7370 -13562 8414 1 OP
rlabel locali -17838 8892 -16746 9030 1 Vdd
rlabel locali -17854 8892 -16746 9030 1 Vdd
rlabel locali -17914 8892 -16746 9216 1 Vdd
rlabel locali -16916 6706 -16882 6842 1 Vss
rlabel metal5 -15198 9332 -15198 9332 1 Vdd
rlabel metal3 -16748 7372 -16660 8416 1 ON
<< end >>
